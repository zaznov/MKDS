module ram_data_gate 
(
input OE, 
input [7:0] IN, 
output [7:0] OUT
);

	assign OUT = (OE ? {8{1'bz}} : IN);
	
endmodule



